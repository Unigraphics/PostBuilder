#################### USER DEFINED EVENTS #####################################
#                                                                            #
#    PURPOSE:                                                                #
#       This file is used in the conversion of post commands contained       #
#       in pre UG V15.0 part files into User Defined Events.                 #
#                                                                            #
##############################################################################


#============================================================================#
#  Created by ling @ Monday, February 22, 2010 6:40:50 PM Pacific Standard Time
#  with Post Builder version 7.5.0.
#============================================================================#


MACHINE FANUC


EVENT auxfun
{
   UI_LABEL "Auxfun"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM auxfun
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Auxfun Value"
   }
   PARAM auxfun_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT clamp
{
   UI_LABEL "Clamp"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM clamp_axis
   {
      TYPE o
      DEFVAL "Xaxis"
      OPTIONS "Xaxis","Yaxis","Zaxis","Aaxis","Baxis","Caxis","Auto"
      UI_LABEL "Clamp Axis"
   }
   PARAM clamp_status
   {
      TYPE o
      DEFVAL "On"
      OPTIONS "On","Off","Axis On","Axis Off"
      UI_LABEL "Clamp Status"
   }
   PARAM clamp_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT coolant
{
   POST_EVENT "coolant_on"
   UI_LABEL "Coolant On"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM coolant_mode
   {
      TYPE o
      DEFVAL "Flood"
      OPTIONS "On","Flood","Mist","Tap","Thru"
      UI_LABEL "Type"
   }
   PARAM coolant_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT coolant_off
{
   UI_LABEL "Coolant Off"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM coolant_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT cutcom
{
   UI_LABEL "Cutter Compensation"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM cutcom_mode
   {
      TYPE o
      DEFVAL "On"
      OPTIONS "Off","On","Left","Right"
      UI_LABEL "Mode"
   }
   PARAM on_option
   {
      TYPE o
      DEFVAL "Before each Engage"
      OPTIONS "Before each Engage","After each Engage","Before 1st Motion"
      UI_LABEL "On"
   }
   PARAM off_option
   {
      TYPE o
      DEFVAL "Before each Retract"
      OPTIONS "Before each Retract","After each Retract","After Last Motion"
      UI_LABEL "Off"
   }
   PARAM Overide_operation_param
   {
      TYPE b
      DEFVAL "TRUE"
      UI_LABEL "Override Operation Parameter"
   }
   PARAM cutcom_adjust_register
   {
      TYPE i
      DEFVAL "0"
      TOGGLE On
      UI_LABEL "Adjust Register"
   }
   PARAM cutcom_plane
   {
      TYPE o
      DEFVAL "NONE"
      OPTIONS "NONE","XY","XZ","YZ"
      UI_LABEL "Plane"
   }
   PARAM full_cutcom_output
   {
      TYPE b
      DEFVAL "FALSE"
      UI_LABEL "Full Cutcom Output"
   }
   PARAM cutcom_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT dnc_header
{
   UI_LABEL "DNC Header"
   CATEGORY MILL DRILL LATHE WEDM
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM dnc_machine_name
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Machine Name"
   }
   PARAM dnc_program_name
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Program Name"
   }
   PARAM dnc_data_type
   {
      TYPE s
      DEFVAL "MPF"
      TOGGLE On
      UI_LABEL "Data Type"
   }
   PARAM dnc_version_number
   {
      TYPE i
      DEFVAL "1"
      TOGGLE On
      UI_LABEL "Version Number"
   }
   PARAM dnc_release_number
   {
      TYPE i
      DEFVAL "1"
      TOGGLE On
      UI_LABEL "Release Number"
   }
   PARAM dnc_user_name
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "User Name"
   }
}


#-----------------------------------------------------------------


EVENT dwell
{
   POST_EVENT "delay"
   UI_LABEL "Dwell"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM delay_mode
   {
      TYPE o
      DEFVAL "Seconds"
      OPTIONS "Seconds","Revolutions"
      UI_LABEL "Dwell Type"
   }
   PARAM delay_value
   {
      TYPE d
      DEFVAL "0.0000"
      UI_LABEL "Dwell Value"
   }
   PARAM delay_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT head
{
   UI_LABEL "Head"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM head_name
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Name"
   }
}


#-----------------------------------------------------------------


EVENT high_speed_setting
{
   UI_LABEL "Sinumerik 840D"
   CATEGORY MILL DRILL
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive"
      UI_LABEL "Status"
   }
   PARAM ude_siemens_tolerance_group
   {
      TYPE g
      DEFVAL "start_closed"
      UI_LABEL "Tolerance"
   }
   PARAM siemens_tol
   {
      TYPE d
      DEFVAL "0.01"
      TOGGLE Off
      UI_LABEL "User Defined Tolerance"
   }
   PARAM ude_siemens_tolerance_group_end
   {
      TYPE g
      DEFVAL "end"
   }
   PARAM ude_siemens_hsm
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "High Speed Machining"
   }
   PARAM siemens_compressor
   {
      TYPE o
      DEFVAL "On"
      OPTIONS "On","Off"
      UI_LABEL "Compressor"
   }
   PARAM siemens_smoothing
   {
      TYPE o
      DEFVAL "On"
      OPTIONS "On","Off"
      UI_LABEL "Smoothing"
   }
   PARAM siemens_feedforward
   {
      TYPE o
      DEFVAL "On"
      OPTIONS "On","Off"
      UI_LABEL "Feed Forward"
   }
   PARAM siemens_5axis_mode
   {
      TYPE o
      DEFVAL "TRAORI"
      OPTIONS "TRAORI","TRAORI2","TRAFOOF","Swiveling"
      UI_LABEL "Transformation"
   }
   PARAM ude_siemens_hsm_end
   {
      TYPE g
      DEFVAL "end"
   }
   PARAM ude_siemens_5axis_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Five Axis Orientation"
   }
   PARAM siemens_ori_coord
   {
      TYPE o
      DEFVAL "Workpiece"
      OPTIONS "Machine","Workpiece"
      UI_LABEL "Coordinate System"
   }
   PARAM siemens_ori_inter
   {
      TYPE o
      DEFVAL "Linear"
      OPTIONS "Linear","Plane"
      UI_LABEL "Interpolation"
   }
   PARAM siemens_ori_def
   {
      TYPE o
      DEFVAL "Rotary Axes"
      OPTIONS "Rotary Axes","Vector"
      UI_LABEL "Definition"
   }
   PARAM siemens_5axis_group_end
   {
      TYPE g
      DEFVAL "end"
   }
   PARAM ude_siemens_feedrate_group
   {
      TYPE g
      DEFVAL "start_closed"
      UI_LABEL "Feed Rate"
   }
   PARAM siemens_feed_definition
   {
      TYPE o
      DEFVAL "Off"
      OPTIONS "On","Off"
      UI_LABEL "Define Feed Rate in Variable"
   }
   PARAM ude_siemens_feedrate_group_end
   {
      TYPE g
      DEFVAL "end"
   }
}


#-----------------------------------------------------------------


EVENT insert
{
   UI_LABEL "Insert"
   PARAM Instruction
   {
      TYPE s
   }
}


#-----------------------------------------------------------------


EVENT instance_operation_handler
{
   UI_LABEL "Instanced Operation Handler"
   PARAM handle_instanced_operations
   {
      TYPE o
      DEFVAL "ON"
      OPTIONS "ON","OFF"
      UI_LABEL "Handle"
   }
}


#-----------------------------------------------------------------


EVENT length_compensation
{
   UI_LABEL "Tool Length Compensation"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM Overide_operation_param
   {
      TYPE b
      DEFVAL "TRUE"
      UI_LABEL "Override Operation Parameter"
   }
   PARAM length_comp_register
   {
      TYPE i
      DEFVAL "2"
      UI_LABEL "Register"
   }
   PARAM length_comp_register_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT lock_axis
{
   UI_LABEL "Lock Axis"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive"
      UI_LABEL "Status"
   }
   PARAM lock_axis
   {
      TYPE o
      DEFVAL "Xaxis"
      OPTIONS "Xaxis","Yaxis","Zaxis","Aaxis","Baxis","Caxis","Fourth","Fifth","Off"
      UI_LABEL "Locked Axis"
   }
   PARAM lock_axis_plane
   {
      TYPE o
      DEFVAL "NONE"
      OPTIONS "XYPLAN","YZPLAN","ZXPLAN","NONE"
      UI_LABEL "Locked Plane"
   }
   PARAM lock_axis_value
   {
      TYPE d
      DEFVAL "0.0000"
      TOGGLE Off
      UI_LABEL "Angle or Coordinate"
   }
}


#-----------------------------------------------------------------


EVENT mill_tool_change
{
   POST_EVENT "load_tool"
   UI_LABEL "Extra Tool Change"
   CATEGORY Mill Drill
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM load_tool_number
   {
      TYPE i
      DEFVAL "0"
      TOGGLE On
      UI_LABEL "Tool Number"
   }
   PARAM tool_z_offset
   {
      TYPE d
      DEFVAL "0.0000"
      TOGGLE Off
      UI_LABEL "Tool Z Offset"
   }
   PARAM tool_adjust_register
   {
      TYPE i
      DEFVAL "0"
      TOGGLE Off
      UI_LABEL "Adjust Register"
   }
   PARAM manual_tool_change
   {
      TYPE b
      DEFVAL "FALSE"
      UI_LABEL "Manual Tool Change"
   }
   PARAM tool_holder
   {
      TYPE i
      DEFVAL "0"
      TOGGLE Off
      UI_LABEL "Holder"
   }
   PARAM tool_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT operator_message
{
   UI_LABEL "Operator Message"
   PARAM operator_message
   {
      TYPE s
      TOGGLE On
      UI_LABEL "Operator Message"
   }
}


#-----------------------------------------------------------------


EVENT opskip_off
{
   UI_LABEL "Optional Skip Off"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM opskip_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT opskip_on
{
   UI_LABEL "Optional Skip On"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM opskip_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT opstop
{
   UI_LABEL "Optional Stop"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM opstop_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT origin
{
   UI_LABEL "Origin"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM X
   {
      TYPE d
      DEFVAL "0.0000"
   }
   PARAM Y
   {
      TYPE d
      DEFVAL "0.0000"
   }
   PARAM Z
   {
      TYPE d
      DEFVAL "0.0000"
   }
   PARAM origin_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT power
{
   UI_LABEL "Power"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM power_value
   {
      TYPE d
      DEFVAL "0.0000"
      UI_LABEL "Power Register"
   }
   PARAM power_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT pprint
{
   UI_LABEL "Pprint"
   PARAM pprint
   {
      TYPE s
      TOGGLE On
      UI_LABEL "Pprint"
   }
}


#-----------------------------------------------------------------


EVENT prefun
{
   UI_LABEL "Prefun"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM prefun
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Prefun Value"
   }
   PARAM prefun_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT program_control
{
   UI_LABEL "Sinumerik Program Control"
   CATEGORY MILL DRILL
   PARAM siemens_program_control
   {
      TYPE b
      DEFVAL "FALSE"
      UI_LABEL "Call External Subroutine for Each Operation"
   }
}


#-----------------------------------------------------------------


EVENT rotate
{
   UI_LABEL "Rotate"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM rotate_axis_type
   {
      TYPE o
      DEFVAL "Table"
      OPTIONS "Table","Head","Aaxis","Baxis","Caxis","Fourth_Axis","Fifth_Axis"
      UI_LABEL "Rotation Axis"
   }
   PARAM rotation_mode
   {
      TYPE o
      DEFVAL "None"
      OPTIONS "None","Angle","Absolute","Incremental"
      UI_LABEL "Type"
   }
   PARAM rotation_direction
   {
      TYPE o
      DEFVAL "CLW"
      OPTIONS "CLW","CCLW","NONE"
      UI_LABEL "Direction"
   }
   PARAM rotation_angle
   {
      TYPE d
      DEFVAL "0.0000"
      TOGGLE On
      UI_LABEL "Angle"
   }
   PARAM rotation_reference_mode
   {
      TYPE b
      DEFVAL "FALSE"
      UI_LABEL "Reference Only - No Output"
   }
   PARAM rotation_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT select_head
{
   UI_LABEL "Select Head"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM head_type
   {
      TYPE o
      DEFVAL "Front"
      OPTIONS "Front","Rear","Right","Left","Side","Saddle"
      UI_LABEL "Head Designation"
   }
   PARAM head_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT sequence_number
{
   UI_LABEL "Sequence Number"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM sequence_mode
   {
      TYPE o
      DEFVAL "N"
      OPTIONS "N","Off","On","Auto"
      UI_LABEL "Number Type"
   }
   PARAM sequence_number
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Number"
   }
   PARAM sequence_increment
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Increment"
   }
   PARAM sequence_frequency
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Frequency"
   }
   PARAM sequence_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT set_axis
{
   UI_LABEL "Set Axis"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM axis_position
   {
      TYPE o
      DEFVAL "ZAXIS"
      OPTIONS "ZAXIS","WAXIS"
      UI_LABEL "Axis"
   }
   PARAM axis_position_value
   {
      TYPE d
      DEFVAL "0.0000"
      TOGGLE On
      UI_LABEL "Position"
   }
}


#-----------------------------------------------------------------


EVENT set_modes
{
   UI_LABEL "Set Modes"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM machine_mode
   {
      TYPE o
      DEFVAL "Mill"
      OPTIONS "Mill","Turn","Punch","Laser","Torch","Wire","Inactive"
      UI_LABEL "Machine Mode"
   }
   PARAM feed_set_mode
   {
      TYPE o
      DEFVAL "Off"
      OPTIONS "Off","IPM","MMPM","IPR","MMPR","FRN","Inactive"
      UI_LABEL "Feed Rate Mode"
   }
   PARAM output_mode
   {
      TYPE o
      DEFVAL "Absolute"
      OPTIONS "Absolute","Increment","Inactive"
      UI_LABEL "Output Mode"
   }
   PARAM arc_mode
   {
      TYPE o
      DEFVAL "Linear"
      OPTIONS "Linear","Circular","Inactive"
      UI_LABEL "Arc Mode"
   }
   PARAM parallel_to_axis
   {
      TYPE o
      DEFVAL "Zaxis"
      OPTIONS "Zaxis","Waxis","Vaxis","Inactive"
      UI_LABEL "Parallel Axis"
   }
   PARAM modes_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT set_polar
{
   UI_LABEL "Set Polar"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM coordinate_output_mode
   {
      TYPE o
      DEFVAL "ON"
      OPTIONS "ON","OFF"
      UI_LABEL "Output Mode"
   }
}


#-----------------------------------------------------------------


EVENT spindle
{
   UI_LABEL "Extra Spindle On"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM spindle_mode
   {
      TYPE o
      DEFVAL "RPM"
      OPTIONS "RPM","SFM","SMM"
      UI_LABEL "Mode"
   }
   PARAM spindle_speed
   {
      TYPE d
      DEFVAL "100.0"
      TOGGLE On
      UI_LABEL "Speed"
   }
   PARAM spindle_maximum_rpm
   {
      TYPE d
      DEFVAL "500.0"
      TOGGLE Off
      UI_LABEL "Maximum Speed"
   }
   PARAM spindle_direction
   {
      TYPE o
      DEFVAL "CLW"
      OPTIONS "CLW","CCLW","NONE"
      UI_LABEL "Direction"
   }
   PARAM spindle_range
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Range"
   }
   PARAM spindle_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT spindle_off
{
   UI_LABEL "Spindle Off"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM spindle_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT stop
{
   UI_LABEL "Stop"
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM stop_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT text
{
   UI_LABEL "User Defined"
   PARAM user_defined_text
   {
      TYPE s
      TOGGLE On
      UI_LABEL "User Defined Command"
   }
}


#-----------------------------------------------------------------


EVENT tool_preselect
{
   UI_LABEL "Tool Preselect"
   CATEGORY MILL DRILL LATHE
   PARAM command_status
   {
      TYPE o
      DEFVAL "Active"
      OPTIONS "Active","Inactive","User Defined"
      UI_LABEL "Status"
   }
   PARAM tool_preselect_number
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Tool Number"
   }
   PARAM tool_preselect_text
   {
      TYPE s
      TOGGLE Off
      UI_LABEL "Text"
   }
}


#-----------------------------------------------------------------


EVENT workpiece_load
{
   UI_LABEL "Load Workpiece"
   CATEGORY MILL DRILL LATHE
   PARAM spindle_number
   {
      TYPE d
      DEFVAL "0.0000"
      TOGGLE OFF
      UI_LABEL "Spindle Number"
   }
}


#-----------------------------------------------------------------


EVENT workpiece_takeover
{
   UI_LABEL "Workpiece Takeover by Spindle 2"
   CATEGORY MILL DRILL LATHE
   PARAM spindle_2_position
   {
      TYPE d
      DEFVAL "0.0000"
      TOGGLE Off
      UI_LABEL "Z Position"
   }
   PARAM takeover_csys
   {
      TYPE o
      DEFVAL "MCS"
      OPTIONS "MCS","MTCS"
      UI_LABEL "Position CSYS"
   }
}


#-----------------------------------------------------------------


EVENT workpiece_unload
{
   UI_LABEL "Unload Workpiece"
   CATEGORY MILL DRILL LATHE
   PARAM spindle_number
   {
      TYPE d
      DEFVAL "0.0000"
      TOGGLE Off
      UI_LABEL "Spindle Number"
   }
}


#-----------------------------------------------------------------


EVENT zero
{
   UI_LABEL "Zero"
   CATEGORY MILL DRILL LATHE
   PARAM work_coordinate_number
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Work Coordinate No."
   }
}


#-----------------------------------------------------------------


SYS_CYCLE Drill_Bore
{
   UI_LABEL "Drill,Bore"
   PARAM ude_siemens_cycle_group
   {
      TYPE g
      DEFVAL "START_OPEN"
      UI_LABEL "Other Parameters"
   }
   PARAM siemens_cycle_rff
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "Retract Feed Rate"
   }
   PARAM ude_siemens_cycle_group_end
   {
      TYPE g
      DEFVAL "end"
   }
}


#-----------------------------------------------------------------


SYS_CYCLE Drill_Bore_Back
{
   UI_LABEL "Drill,Bore,Back"
   PARAM ude_siemens_cycle_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Retract Distance"
   }
   PARAM siemens_cycle_rpa
   {
      TYPE d
      DEFVAL "0.0"
      UI_LABEL "X"
   }
   PARAM siemens_cycle_rpo
   {
      TYPE d
      DEFVAL "0.0"
      UI_LABEL "Y"
   }
   PARAM siemens_cycle_rpap
   {
      TYPE d
      DEFVAL "0.0"
      UI_LABEL "Z"
   }
   PARAM ude_siemens_cycle_group_end
   {
      TYPE g
      DEFVAL "end"
   }
}


#-----------------------------------------------------------------


SYS_CYCLE Drill_Bore_Nodrag
{
   UI_LABEL "Drill,Bore,Nodrag"
   PARAM ude_siemens_cycle_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Retract Distance"
   }
   PARAM siemens_cycle_rpa
   {
      TYPE d
      DEFVAL "0.0"
      UI_LABEL "X"
   }
   PARAM siemens_cycle_rpo
   {
      TYPE d
      DEFVAL "0.0"
      UI_LABEL "Y"
   }
   PARAM siemens_cycle_rpap
   {
      TYPE d
      DEFVAL "0.0"
      UI_LABEL "Z"
   }
   PARAM ude_siemens_cycle_group_end
   {
      TYPE g
      DEFVAL "end"
   }
}


#-----------------------------------------------------------------


SYS_CYCLE Drill_Deep
{
   UI_LABEL "Drill,Deep"
   PARAM ude_siemens_cycle_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Other Parameters"
   }
   PARAM siemens_cycle_dts_mode
   {
      TYPE o
      DEFVAL "Off"
      OPTIONS "Off","On","Seconds","Revolutions"
      UI_LABEL "Top Dwell"
   }
   PARAM siemens_cycle_dts
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Top Dwell Value"
   }
   PARAM siemens_cycle_o_dtd_mode
   {
      TYPE o
      DEFVAL "Off"
      OPTIONS "Off","On","Seconds","Revolutions"
      UI_LABEL "Final Dwell"
   }
   PARAM siemens_cycle_o_dtd
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Final Dwell Value"
   }
   PARAM siemens_cycle_frf
   {
      TYPE d
      DEFVAL "1"
      UI_LABEL "Feed Rate Factor"
   }
   PARAM siemens_cycle_o_dis1
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "Step Clearance"
   }
   PARAM ude_siemens_cycle_group_end
   {
      TYPE g
      DEFVAL "end"
   }
}


#-----------------------------------------------------------------


SYS_CYCLE Drill_Deep_Breakchip
{
   UI_LABEL "Drill,Deep,BreakChip"
   PARAM ude_siemens_cycle_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Other Parameters"
   }
   PARAM siemens_cycle_o_dtd_mode
   {
      TYPE o
      DEFVAL "Off"
      OPTIONS "Off","On","Seconds","Revolutions"
      UI_LABEL "Final Dwell"
   }
   PARAM siemens_cycle_o_dtd
   {
      TYPE i
      DEFVAL "0"
      UI_LABEL "Final Dwell Value"
   }
   PARAM siemens_cycle_frf
   {
      TYPE d
      DEFVAL "1"
      UI_LABEL "Feed Rate Factor"
   }
   PARAM siemens_cycle_o_vrt
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "Step Retract Value"
   }
   PARAM ude_siemens_cycle_group_end
   {
      TYPE g
      DEFVAL "end"
   }
}


#-----------------------------------------------------------------


SYS_CYCLE Drill_Tap
{
   UI_LABEL "Drill,Tap"
   PARAM ude_siemens_thread_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Pitch"
   }
   PARAM siemens_cycle_mpit
   {
      TYPE i
      DEFVAL "3"
      TOGGLE Off
      UI_LABEL "Thread Size"
   }
   PARAM siemens_cycle_o_ptab
   {
      TYPE o
      DEFVAL "Post Defined"
      OPTIONS "Post Defined","Millimeter","Groove per Inch","Inch per Revolution"
      UI_LABEL "Pitch"
   }
   PARAM siemens_cycle_pit
   {
      TYPE d
      DEFVAL "0.0"
      UI_LABEL "Pitch Value"
   }
   PARAM ude_siemens_thread_group_end
   {
      TYPE g
      DEFVAL "end"
   }
   PARAM ude_siemens_float_group
   {
      TYPE g
      DEFVAL "start_closed"
      UI_LABEL "Float Tap Parameters"
   }
   PARAM siemens_cycle_sdr
   {
      TYPE o
      DEFVAL "Reversal"
      OPTIONS "CLW","CCLW","Reversal"
      UI_LABEL "Spindle Retract Direction"
   }
   PARAM siemens_cycle_enc
   {
      TYPE o
      DEFVAL "Use Encoder-Dwell Off"
      OPTIONS "Use Encoder-Dwell Off","Use Encoder-Dwell On","No Encoder-Feed Rate before Cycle","No Encoder-Feed Rate in Cycle"
      UI_LABEL "Encoder"
   }
   PARAM ude_siemens_float_group_end
   {
      TYPE g
      DEFVAL "end"
   }
   PARAM ude_siemens_rigid_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Rigid Tap Parameters"
   }
   PARAM siemens_cycle_o_var1
   {
      TYPE o
      DEFVAL "Single Pass"
      OPTIONS "Single Pass","Break Chip","Remove Chip"
      UI_LABEL "Type"
   }
   PARAM siemens_cycle_poss
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "Spindle Orient Angle"
   }
   PARAM siemens_cycle_sst1
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "Spindle Retract Speed"
   }
   PARAM siemens_cycle_o_dam
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "Deep Hole Incremental Depth"
   }
   PARAM siemens_cycle_o_vrt
   {
      TYPE d
      DEFVAL "0.0"
      TOGGLE Off
      UI_LABEL "Break Chip Retract Value"
   }
   PARAM ude_siemens_rigid_group_end
   {
      TYPE g
      DEFVAL "end"
   }
   PARAM ude_siemens_other_group
   {
      TYPE g
      DEFVAL "start_open"
      UI_LABEL "Other Parameters"
   }
   PARAM siemens_cycle_sdac
   {
      TYPE o
      DEFVAL "CLW"
      OPTIONS "CLW","CCLW","Off"
      UI_LABEL "Spindle Direction After Cycle"
   }
   PARAM siemens_cycle_o_techno
   {
      TYPE i
      DEFVAL "0"
      TOGGLE Off
      UI_LABEL "Technological Setting"
   }
   PARAM ude_siemens_other_end
   {
      TYPE g
      DEFVAL "end"
   }
}


#-----------------------------------------------------------------


