#############################################################################################
#
#	Copyright 2014-2019 Siemens Product Lifecycle Management Software Inc.
#				All Rights Reserved.
#
#############################################################################################

MACHINE GENERIC
