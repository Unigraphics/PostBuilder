#############################################################################################
#
#	Customer Data
#
#	Company         :
#	Address         :
#	Contact person  :
#	Phone           :
#	Fax             :
#	Mail            :
#
#############################################################################################
#
#	Copyright 2014-2019 Siemens Product Lifecycle Management Software Inc.
#				All Rights Reserved.
#
#############################################################################################

MACHINE Default
